import("net/tBuffer.cdl");
import("netinet/tNetworkTimer.cdl");

import("netdev/if_mbed/tIfMbed.cdl");
import("netdev/if_mbed/tIfMbedAdapter.cdl");
import("net/tEthernet.cdl");
import("netinet/tArp.cdl");

cell tKernel Kernel {
};

/**
*   イーサネット層
*
**/

[allocator(eArpInput.arpInput.inputp=NetworkBuffer.eNetworkAlloc,
           eArpOutput.arpResolve.outputp=NetworkBuffer.eNetworkAlloc)]
cell tArp Arp {

    cEthernetRawOutput = EthernetOutputTaskBody.eRawOutput;
    //cIPv4Functions = IPv4Functions.eFunctions;

    cNetworkTimer = NetworkTimer.eNetworkTimer[1];
    cArpSemaphore = ArpSemaphore.eSemaphore;

    arpEntry = 10;
};

cell tTask EthernetInputTask {

    cTaskBody = EthernetInputTaskBody.eTaskBody;

    attribute = C_EXP("TA_HLNG|TA_ACT");
    priority  = C_EXP("ETHER_INPUT_PRIORITY");
    stackSize = C_EXP("ETHER_INPUT_STACK_SIZE");
};

cell tEthernetInputTaskBody EthernetInputTaskBody {

    cTaskNetworkTimer = NetworkTimerTask.eTask;
    cTaskEthernetOutput = EthernetOutputTask.eTask;
    cSemaphoreReceive = SemaphoreNicReceive.eSemaphore;
    cNicDriver = IfMbed.eNicDriver;

    cArpInput = Arp.eArpInput;
    //cIPv4Input = IPv4Input.eIPv4Input;
};

cell tTask EthernetOutputTask {

    cTaskBody = EthernetOutputTaskBody.eTaskBody;

    attribute = C_EXP("TA_HLNG");
    priority  = C_EXP("ETHER_OUTPUT_PRIORITY");
    stackSize = C_EXP("ETHER_OUTPUT_STACK_SIZE");
};

[allocator(eRawOutput.ethernetRawOutput.outputp=NetworkBuffer.eNetworkAlloc)]
cell tEthernetOutputTaskBody EthernetOutputTaskBody {

    cNicDriver = IfMbed.eNicDriver;
    cSemaphoreSend = SemaphoreNicSend.eSemaphore;
    cSemaphoreTcppost = SemaphoreTcppost.eSemaphore;
    cDataqueue = DataqueueEthernet.eDataqueue;
};

//[allocator(eEthernetOutput.ethernetOutput.outputp=NetworkBuffer.eNetworkAlloc)]
cell tEthernetOutput EthernetOutput {

    cNicDriver = IfMbed.eNicDriver;
    cArpOutput = Arp.eArpOutput;
    cRawOutput = EthernetOutputTaskBody.eRawOutput;
};

/**
*   物理層
*   tNetworkInterfaceContllor (tIfMbed)
**/

[allocator(eNicDriver.start.outputp=NetworkBuffer.eNetworkAlloc,
			eNicDriver.read.inputp=NetworkBuffer.eNetworkAlloc)]
cell tIfMbed IfMbed {

	cSemaphoreSend 		= SemaphoreNicSend.eSemaphore;
	//ciSemaphoreReceive 	= SemaphoreNicReceive.eiSemaphore;
	cSemaphoreReceive 	= SemaphoreNicReceive.eSemaphore;
	cInterruptRequest 	= NicInterrupt.eInterruptRequest;

    cNetworkTimer = NetworkTimer.eNetworkTimer[0];

    cTask = IfMbedPhyTask.eTask;
};

cell tTask IfMbedPhyTask {

    cTaskBody = IfMbedPhyTaskBody.eTaskBody;

    attribute = C_EXP("TA_NULL");
    priority  = C_EXP("IF_MBED_PHY_PRIORITY");
    stackSize = C_EXP("IF_MBED_PHY_STACK_SIZE");
};

cell tIfMbedPhyTaskBody IfMbedPhyTaskBody {
};

cell tIfMbedAdapter IfMbedAdapter {

	cNicDriver = IfMbed.eNicDriver;
};

/*
*   Dataquque, Semaphore etc.
*/
cell tSemaphore ArpSemaphore{
    attribute       = C_EXP("TA_TPRI");
    initialCount    = 1;
    maxCount        = 1;
};
cell tDataqueue DataqueueEthernet{

    attribute                   = C_EXP("TA_NULL");
    dataCount                   = 1;
    dataqueueManagementBuffer   = C_EXP("NULL");
};
cell tSemaphore SemaphoreNicSend {

    attribute 		= C_EXP("TA_TPRI");
    initialCount 	= 1;
    maxCount 		= 1;
};
cell tSemaphore SemaphoreNicReceive {

    attribute 		= C_EXP("TA_TPRI");
    initialCount 	= 0;
    maxCount 		= 1;
};
cell tSemaphore SemaphoreTcppost {

    attribute       = C_EXP("TA_TPRI");
    initialCount    = 0;
    maxCount        = 1;
};
cell tISRWithInterruptRequest NicInterrupt {

	ciISRBody = IfMbed.eiBody;

	interruptNumber 	= (0x200);
	interruptAttribute 	= C_EXP("TA_ENAINT");
	interruptPriority 	= -8;
};

/**
*   タイマ組み上げ宣言
**/
cell tNetworkTimer NetworkTimer{
    //cTCPTask = TCPTask.eTask;

    /* 有効なネットワークタイマ宣言 */
    cCallTimerFunction[0] = IfMbed.eWatchdogTimer;
    cCallTimerFunction[1] = Arp.eArpTimer;
    //cCallTimerFunction[2] = IPv4RoutingTable.eRoutingTableTimer;
    //cCallTimerFunction[3] = TCPOutputBody.eCallTimerFunction;

    cSemaphoreNetworkTimer  = SemaphoreNetworkTimer.eSemaphore;
    ciSemaphoreNetworkTimer = SemaphoreNetworkTimer.eiSemaphore;
    cSemaphoreCalloutLock   = SemaphoreCalloutLock.eSemaphore;
};
