import_C("netinet/tecs_if_ether.h");

celltype tArp {

    //call sIPv4Functions cIPv4Functions;
    call sEthernetRawOutput cEthernetRawOutput;

    //call sNetworkTimer cNetworkTimer;
    call sSemaphore cArpSemaphore;

    entry sArpInput eArpInput;
    entry sArpOutput eArpOutput;
    //entry sCallTimerFunction eArpTimer;

    attr{
        int32_t arpEntry;
    };

    var{
        [size_is(arpEntry)]T_ARP_ENTRY *arp_cache;
    };
};