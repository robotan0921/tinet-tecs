import_C("net/tecs_net.h");

import("net/tBuffer.cdl");
import("netinet/tNetworkTimer.cdl");

import("netdev/if_mbed/tIfMbed.cdl");
import("netdev/if_mbed/tIfMbedAdapter.cdl");

import("net/tEthernet.cdl");

import("netinet/tIPv4.cdl");
import("netinet/tArp.cdl");
import("netinet/tIPv4InputAdapter.cdl");

import("netinet/tTCP.cdl");

//TCPCEPの数
const uint32_t NUM_TCPCEP = 1;

cell tKernel Kernel {
};

/**
*   トランスポート層
*
**/
[allocator(eInput.TCPInput.inputp=NetworkBuffer.eNetworkAlloc),generate(RepeatPlugin ,"count = NUM_TCPCEP")] //TODO: 逆リクワイアsendが使えないためとりあえず
cell tTCPInput TCPInput {

    //cCEPInput[0]  = TCPCEP_000.eInput;
    cIPv4CheckSum = IPv4Functions.eCheckSum;
    cTCPRespond   = TCPOutputBody.eTCPOutput;
};

[generate(RepeatPlugin ,"count = NUM_TCPCEP"),allocator(eTCPOutput.output.outputp=NetworkBuffer.eNetworkAlloc,
                                                        eTCPOutput.respond.outputp=NetworkBuffer.eNetworkAlloc)]
cell tTCPOutputBody TCPOutputBody {
    //cTCPOutputStart[0] = TCPCEP_000.eTCPOutputStart;
    cIPv4Output        = IPv4Output.eOutput;
    cIPv4CheckSum      = IPv4Functions.eCheckSum;
    cSemaphore         = SemaphoreTcppost.eSemaphore;
    cNetworkTimer      = NetworkTimer.eNetworkTimer[3];
    cTCPFunctions      = TCPFunctions.eTCPFunctions;
};

cell tTask TCPTask {

    cTaskBody = TCPOutputBody.eTaskBody;

    attribute = C_EXP("TA_NULL");
    priority  = 5;
    stackSize = 1024;
};

cell tTCPFunctions TCPFunctions {
};

/**
*   ネットワーク層
*
**/
const T_IN4_ADDR MYIP4ADDRESS = C_EXP("MAKE_IPV4_ADDR(192,168,1,200)");
const T_IN4_ADDR MYIP4MASK    = C_EXP("MAKE_IPV4_ADDR(255,255,255,0)");
const T_IN4_ADDR MYIP4GATAWAY = C_EXP("MAKE_IPV4_ADDR(192,168,1,1)");

cell tIPv4RoutingTable IPv4RoutingTable {

    cSemaphore    = SemaphoreIPv4Routing.eSemaphore;
    cNetworkTimer = NetworkTimer.eNetworkTimer[2];

    numStaticEntry   = 3;
    numRedirectEntry = 1;
    timeout          = 10;
    staticRoutingTable = {
        {0, 0, C_EXP("MYIP4GATAWAY"), 0, C_EXP("IN_RTF_DEFINED")},
        {C_EXP("MYIP4ADDRESS &MYIP4MASK"), C_EXP("MYIP4MASK"), 0, 0, C_EXP("IN_RTF_DEFINED")},
        {C_EXP("0xffffffff,0xffffffff,0"), 0, C_EXP("IN_RTF_DEFINED")}
    };
};

cell tIPv4Functions IPv4Functions {

    IPv4AddressInit = MYIP4ADDRESS;
    IPv4MaskInit    = MYIP4MASK;
    IPv4GatawayInit = MYIP4GATAWAY;
};

[allocator(eICMP4.input.inputp=NetworkBuffer.eNetworkAlloc,
           eICMP4Error.error.inputp=NetworkBuffer.eNetworkAlloc)]
cell tICMP4 ICMP4 {

    //cTCPInput      = TCPInput.eInput;
    cIPv4Reply     = IPv4Output.eOutput;
    cIPv4Functions = IPv4Functions.eFunctions;
};

[allocator(eIPv4Input.IPv4Input.inputp=NetworkBuffer.eNetworkAlloc)]
cell tIPv4Input IPv4Input {

    cFunctions  = IPv4Functions.eFunctions;
    cICMP4      = ICMP4.eICMP4;
    cICMP4Error = ICMP4.eICMP4Error;
    //cUDPInput   = UDPInput.eInput;
    //cTCPInput   = TCPInput.eInput;
};

[allocator(eOutput.IPv4Output.outputp=NetworkBuffer.eNetworkAlloc,
           eOutput.IPv4Reply.outputp=NetworkBuffer.eNetworkAlloc)]
cell tIPv4Output IPv4Output {

    cEthernetOutput = EthernetOutput.eEthernetOutput;
    cFunctions      = IPv4Functions.eFunctions;
    cRoutingTable   = IPv4RoutingTable.eRoutingTable;
    cIPv4CheckSum   = IPv4Functions.eCheckSum;
};

/**
*   イーサネット層
*
**/

[allocator(eArpInput.arpInput.inputp=NetworkBuffer.eNetworkAlloc,
           eArpOutput.arpResolve.outputp=NetworkBuffer.eNetworkAlloc)]
cell tArp Arp {

    cEthernetRawOutput = EthernetOutputTaskBody.eRawOutput;
    cFunctions = IPv4Functions.eFunctions;

    cNetworkTimer = NetworkTimer.eNetworkTimer[1];
    cArpSemaphore = ArpSemaphore.eSemaphore;

    arpEntry = 10;
};

cell tTask EthernetInputTask {

    cTaskBody = EthernetInputTaskBody.eTaskBody;

    attribute = C_EXP("TA_HLNG|TA_ACT");
    priority  = C_EXP("ETHER_INPUT_PRIORITY");
    stackSize = C_EXP("ETHER_INPUT_STACK_SIZE");
};

cell tEthernetInputTaskBody EthernetInputTaskBody {

    cTaskNetworkTimer = NetworkTimerTask.eTask;
    cTaskEthernetOutput = EthernetOutputTask.eTask;
    cSemaphoreReceive = SemaphoreNicReceive.eSemaphore;
    cNicDriver = IfMbed.eNicDriver;

    cArpInput = Arp.eArpInput;
    cIPv4Input = IPv4Input.eIPv4Input;
};

cell tTask EthernetOutputTask {

    cTaskBody = EthernetOutputTaskBody.eTaskBody;

    attribute = C_EXP("TA_HLNG");
    priority  = C_EXP("ETHER_OUTPUT_PRIORITY");
    stackSize = C_EXP("ETHER_OUTPUT_STACK_SIZE");
};

[allocator(eRawOutput.ethernetRawOutput.outputp=NetworkBuffer.eNetworkAlloc)]
cell tEthernetOutputTaskBody EthernetOutputTaskBody {

    cNicDriver = IfMbed.eNicDriver;
    cSemaphoreSend = SemaphoreNicSend.eSemaphore;
    cSemaphoreTcppost = SemaphoreTcppost.eSemaphore;
    cDataqueue = DataqueueEthernet.eDataqueue;
};

[allocator(eEthernetOutput.ethernetOutput.outputp=NetworkBuffer.eNetworkAlloc)]
cell tEthernetOutput EthernetOutput {

    cNicDriver = IfMbed.eNicDriver;
    cArpOutput = Arp.eArpOutput;
    cRawOutput = EthernetOutputTaskBody.eRawOutput;
};

/**
*   物理層
*   tNetworkInterfaceContllor (tIfMbed)
**/

[allocator(eNicDriver.start.outputp=NetworkBuffer.eNetworkAlloc,
			eNicDriver.read.inputp=NetworkBuffer.eNetworkAlloc)]
cell tIfMbed IfMbed {

	ciSemaphoreSend 	= SemaphoreNicSend.eiSemaphore;
	cSemaphoreReceive 	= SemaphoreNicReceive.eSemaphore;
	cInterruptRequest 	= NicInterrupt.eInterruptRequest;

    cNetworkTimer = NetworkTimer.eNetworkTimer[0];

    cTask = IfMbedPhyTask.eTask;
};

cell tTask IfMbedPhyTask {

    cTaskBody = IfMbedPhyTaskBody.eTaskBody;

    attribute = C_EXP("TA_NULL");
    priority  = C_EXP("IF_MBED_PHY_PRIORITY");
    stackSize = C_EXP("IF_MBED_PHY_STACK_SIZE");
};

cell tIfMbedPhyTaskBody IfMbedPhyTaskBody {
};


/*
*   Adapters
*/
cell tIfMbedAdapter IfMbedAdapter {

	cNicDriver = IfMbed.eNicDriver;
};
cell tIPv4InputAdapter IPv4InputAdapter {

    cIPv4Input = IPv4Input.eIPv4Input;
};
/*
*   Dataquque, Semaphore etc.
*/
cell tSemaphore SemaphoreTcppost {

    attribute       = C_EXP("TA_TPRI");
    initialCount    = 0;
    maxCount        = 1;
};
cell tSemaphore SemaphoreIPv4Routing {

    attribute       = C_EXP("TA_TPRI");
    initialCount    = 1;
    maxCount        = 1;
};
cell tSemaphore ArpSemaphore {

    attribute       = C_EXP("TA_TPRI");
    initialCount    = 1;
    maxCount        = 1;
};
cell tDataqueue DataqueueEthernet{

    attribute                   = C_EXP("TA_NULL");
    dataCount                   = 1;
    dataqueueManagementBuffer   = C_EXP("NULL");
};
cell tSemaphore SemaphoreNicSend {

    attribute 		= C_EXP("TA_TPRI");
    initialCount 	= 1;
    maxCount 		= 1;
};
cell tSemaphore SemaphoreNicReceive {

    attribute 		= C_EXP("TA_TPRI");
    initialCount 	= 0;
    maxCount 		= 1;
};
cell tISRWithInterruptRequest NicInterrupt {

	ciISRBody = IfMbed.eiBody;

	interruptNumber 	= (0x200);
	interruptAttribute 	= C_EXP("TA_ENAINT");
	interruptPriority 	= -8;
};

/**
*   タイマ組み上げ宣言
**/
cell tNetworkTimer NetworkTimer{
    cTCPTask = TCPTask.eTask;

    /* 有効なネットワークタイマ宣言 */
    cCallTimerFunction[0] = IfMbed.eWatchdogTimer;
    cCallTimerFunction[1] = Arp.eArpTimer;
    cCallTimerFunction[2] = IPv4RoutingTable.eRoutingTableTimer;
    cCallTimerFunction[3] = TCPOutputBody.eCallTimerFunction;

    cSemaphoreNetworkTimer  = SemaphoreNetworkTimer.eSemaphore;
    ciSemaphoreNetworkTimer = SemaphoreNetworkTimer.eiSemaphore;
    cSemaphoreCalloutLock   = SemaphoreCalloutLock.eSemaphore;
};
